module cpu (
    input logic clk,
    input logic reset
);


endmodule
